module mod

pub fn mod_fun() {}
