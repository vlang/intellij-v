module main

struct Foo {}
interface Ifoo {}
union Ufoo {}
enum Efoo {}

struct f {}
interface i {}
union u {}
enum e {}
