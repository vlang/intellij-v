module second

import first

pub fn util() {
	first.util()
}
