module main

type <error descr="Type alias name must start with uppercase letter">mystring</error> = string
