module namingConventions

const named_constant = 100
const ok_constant = 100
