module main
fn main() {
    <error descr="Variable name cannot contain uppercase letters, use snake_case instead">InvalidVarName</error> := 1
}