module stubs

pub struct UnknownCDeclaration {
pub mut:
	unknown_field &UnknownCDeclaration
}

pub fn (c &UnknownCDeclaration) unknown_method()
