module inner

pub fn inner() {
	println!("inner");
}
