module parser

fn main() {
	`0`
	`\0`
	`\``
	`\n`
	`\a`
	`🚀`

	`\x61`
	`\141`
	`\u0061`

	`\u2605`
	`\u2605`
	`\xe2\x98\x85`
	`\342\230\205`
	`\uFFFF`
}
