module builtin

fn println(s string) {}
