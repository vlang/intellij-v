module inner

pub struct Foo {

}

pub fn (a []Foo) foo() {

}

pub fn (a map[string]Foo) boo() {

}
