module annotators

enum <warning descr="Enum must have at least one field">Empty</warning> {}

enum WithFields {
	red
	green
}
