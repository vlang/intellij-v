module main

enum Colors {
	red
	green
}
fn main() {
	mut color := Colors.red
	expr_type(color, 'Colors')
}
