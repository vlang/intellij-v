module postfix

names := [1, 2, 3]

for name in names {
	<caret>
}
