module simple

pub struct SimpleStruct {

}

pub fn simple_func() {}
