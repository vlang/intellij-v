module main

fn main() {
	$for field in fields {

	}

	$for i := 0; i < 100; i++ {

	}

	$for i, key in value {

	}
}
