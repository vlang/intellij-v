module parser

struct Foo {}

fn main() {
	for i := 0; i < 100; {
		Foo{}
	}
}
