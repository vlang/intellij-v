module mymodule

pub fn my_func() {
	return 42
}
