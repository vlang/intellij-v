module main

fn pascal_case() {}
fn camel_case() {}
fn snake_case() {}
fn invalid_snake_case() {}
