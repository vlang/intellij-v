module annotators

struct Foo {
pub mut:
	a int
pub mut:
	b int
}
