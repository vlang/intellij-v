module main

fn pascal_case() {}
fn camel_case() {}
fn snake_case() {}
fn invalid_snake_case() {}

fn (s string) pascal_case() {}
fn (s string) camel_case() {}
fn (s string) snake_case() {}
fn (s string) invalid_snake_case() {}
