module mod
