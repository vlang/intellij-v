module namingConventions

fn C.foo() {}
fn JS.foo() {}
fn WASM.foo() {}

struct C.Name {}
struct JS.Name {}
struct WASM.Name {}

type C.void = void
