module with_src

fn with_src_func() {}
