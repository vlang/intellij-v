module main

fn main() {
	unsafe {
		println(nil)
	}
}
