module main

type Mystring = string
