module main

type Keyword = int

fn import() {}
fn struct() {}
fn implements() {}
fn union() {}
fn interface() {}
fn enum() {}
fn const() {}
fn type() {}
fn fn() {}
fn return() {}
fn select() {}
fn match() {}
fn or() {}
fn if() {}
fn else() {}
fn goto() {}
fn assert() {}
fn for() {}
fn break() {}
fn continue() {}
fn unsafe() {}
fn defer() {}
fn go() {}
fn spawn() {}
fn rlock() {}
fn lock() {}
fn as() {}
fn in() {}
fn is() {}
fn nil() {}
fn none() {}
fn static() {}
fn shared() {}
fn atomic() {}
fn dump() {}
fn sizeof() {}
fn typeof() {}
fn isreftype() {}
fn module() {}
fn true() {}
fn false() {}
fn pub() {}
fn mut() {}
fn volatile() {}
// fn asm() {}
// fn __global() {}
// fn __offsetof() {}

fn (k Keyword) import() {}
fn (k Keyword) struct() {}
fn (k Keyword) implements() {}
fn (k Keyword) union() {}
fn (k Keyword) interface() {}
fn (k Keyword) enum() {}
fn (k Keyword) const() {}
fn (k Keyword) type() {}
fn (k Keyword) fn() {}
fn (k Keyword) return() {}
fn (k Keyword) select() {}
fn (k Keyword) match() {}
fn (k Keyword) or() {}
fn (k Keyword) if() {}
fn (k Keyword) else() {}
fn (k Keyword) goto() {}
fn (k Keyword) assert() {}
fn (k Keyword) for() {}
fn (k Keyword) break() {}
fn (k Keyword) continue() {}
fn (k Keyword) unsafe() {}
fn (k Keyword) defer() {}
fn (k Keyword) go() {}
fn (k Keyword) spawn() {}
fn (k Keyword) rlock() {}
fn (k Keyword) lock() {}
fn (k Keyword) as() {}
fn (k Keyword) in() {}
fn (k Keyword) is() {}
fn (k Keyword) nil() {}
fn (k Keyword) none() {}
fn (k Keyword) static() {}
fn (k Keyword) shared() {}
fn (k Keyword) atomic() {}
fn (k Keyword) dump() {}
fn (k Keyword) sizeof() {}
fn (k Keyword) typeof() {}
fn (k Keyword) isreftype() {}
fn (k Keyword) module() {}
fn (k Keyword) true() {}
fn (k Keyword) false() {}
fn (k Keyword) pub() {}
fn (k Keyword) mut() {}
fn (k Keyword) volatile() {}
// fn (k Keyword) asm() {}
// fn __global() {}
// fn __offsetof() {}