module mymodule2

pub fn my_func2() {
	return 42
}
