module builtin

interface IError {}
