module builtin

pub struct string {

}
