module main

struct Test {
pub:
	name string
}

fn main() {
	match 100 {
		200 {}
	}

	test := Test{
		name: ''
	}
}
