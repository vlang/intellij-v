module postfix

name_to_id := map[string]int{}

for key, id in name_to_id {
	<caret>
}
