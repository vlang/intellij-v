module postfix

mp := map[string]int{}

for key, value in mp {
	<caret>
}