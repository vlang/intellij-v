module main

import os
import os as os2

import v.doc
import v.doc as vdoc

fn main() {
	os.args
	os2.args

	doc.Doc{}
	vdoc.Doc{}
}
