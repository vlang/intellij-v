module main

import /*caret*/mod

mod.mod_fun()
