module builtin

pub fn println(s string) {}
