module annotators

mp := map[string]int{}

for _, value in mp {

}

for key, value in mp {

}