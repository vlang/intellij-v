module main

struct Test {
	name string
	name string
	name string
}

enum Colors {
	red
	blue
	ye_l_llow
	blue
}
