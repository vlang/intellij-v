module types

a := 100
expr_type(a++, 'int')
