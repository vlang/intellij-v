module postfix

name_to_id := map[string]int{}

name_to_id.for<caret>
