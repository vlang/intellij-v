module postfix

names := [1, 2, 3]

names.for<caret>
