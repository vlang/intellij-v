module main

fn main() {
	if i in [
		Test{
			text_document: doc_id
		},
		Test{
			text_document: doc_id
		},
	] {
	}

	if _ := code_lens(Test{ text_document: doc_id }, mut writer) {
		println('')
	} else {
		println('')
	}

	for i := 0; i < 100; i++ {
		idxs << RepIndex{
			idx: idx
			val_idx: rep_i
		}
	}

	match '' {
		'array' {
			idxs << RepIndex{
				idx: idx
				val_idx: rep_i
			}
		}
		else {}
	}

	fun(if v { 1 } else { 0 })
}
