module postfix

arr := [1, 2, 3]

arr.for<caret>
