module nested

pub fn nested_fn() {
	println("nested_fun");
}
