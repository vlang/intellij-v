module types

fn main() {
	expr_type(chan int{}, 'chan int')
}
