module postfix

mp := map[string]int{}

mp.for<caret>
