module types

expr_type(_likely_(a > 100), 'bool')
expr_type(_unlikely_(a > 100), 'bool')
