module simple

pub fn simple_func() {}
