module new

a := 100

dump(100)
dump(a + 100)
