module main

struct Foo {}
interface Ifoo {}
union Ufoo {}
enum Efoo {
	red
}

struct f {}
interface i {}
union u {}
enum e {
	red
}
