module namingConventions

const <error descr="Constant name cannot contain uppercase letters, use snake_case instead">NamedConstant</error> = 100
const ok_constant = 100
