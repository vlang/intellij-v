module json
