module sub

pub fn sub() {
	println!("sub");
}
