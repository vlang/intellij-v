module namingConventions

fn C.foo() {}
fn JS.foo() {}

struct C.Name {}
struct JS.Name {}

type C.void = void
