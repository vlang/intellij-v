module validity

mut arr := []int{}
arr << 1

mut arr_mut := []int{}
arr_mut << 1
