module new

import gx

fn main() {
	if book is fn () {
	}
	if book == Book{} {
	}
	if book is Book {
	}
	if author == name {
		hello := 100
	}
	name := 100
	match name {
		Book {
			println()
		}
		Book, Book {}
		else {}
	}

	match kind {
		.points {
			return gx.TextCfg{}
		}
		.moves {
			return gx.TextCfg{}
		}
	}

	possible_moves := [1, 2, 3]
	for move_idx in 0 .. possible_moves.len {
		1
	}

	write8(match true {
		size == 1 && is_signed { 0xbe }
		else { 0x8b }
	})

	match {
		'name': 100
	} {
		map[string]int {}
		fn () {}
		else {}
	}
	match Book {
		map[string]int {}
	}
	a := {
		'name': 100
	}
}

