module first

import second

pub fn util() {
	second.util()
}
