module parser

struct User {}

fn User.new() User {
	return User{}
}

user := User.new()