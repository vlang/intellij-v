module types

fn main() {
	for i in 0 .. 100 {
		expr_type(i, 'int')
	}
}
