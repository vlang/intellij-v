module sub

struct Sub {

}
