module postfix

arr := [1, 2, 3]

for value in arr {
	<caret>
}