module stubs

pub struct UnknownCDeclaration {
pub:
	unknown_field &UnknownCDeclaration
}

pub fn (c &UnknownCDeclaration) unknown_method()
